library verilog;
use verilog.vl_types.all;
entity busloko is
end busloko;
