class sequence extends uvm_sequence;

endclass : sequence