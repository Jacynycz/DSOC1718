library verilog;
use verilog.vl_types.all;
entity bfm_sv_unit is
end bfm_sv_unit;
