library verilog;
use verilog.vl_types.all;
entity tester_sv_unit is
end tester_sv_unit;
