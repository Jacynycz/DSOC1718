`include "uvm_macros.sv"
package my_package;
import uvm_pkg::*;
`include "general_seq_item.sv"
`include "add_seq_item.sv"
`include "and_seq_item.sv"
`include "xor_seq_item.sv"
`include "mul_seq_item.sv"
endpackage 