library verilog;
use verilog.vl_types.all;
entity coverage_sv_unit is
end coverage_sv_unit;
