
package imports;
	parameter version = "1.0";
	// Sequence items
	`include "general_seq_item.sv"
	`include "add_seq_item.sv"
	`include "xor_seq_item.sv"
	`include "mul_seq_item.sv"
	`include "and_seq_item.sv"
	
	// driver


	// monitors


	// scoreboard


	// agent


endpackage