`include "uvm_macros.svh"
module top;
import uvm_pkg::*;
import my_package::*;

initial
begin
	
end
endmodule