
package imports;
	parameter version = "1.0";
	`include "transaction.sv"
	`include "driver.sv"
endpackage